module encoder_4x2(d0,d1,d2,d3,q0,q1);
  input d0,d1,d2,d3;
  output q0,q1;
  assign q0 = d3|d1;
  assign q1 = d3|d2;
endmodule
