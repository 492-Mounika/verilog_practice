module counter(
    input wire clk,
    input wire reset,
    input wire valid,
    output reg [3:0]count
);
always @(posedge clk) begin
    if (reset) begin
        count <= 4'b0000;
    end
    else begin
        if (valid) begin
            count <= count+1;
        end
    end
end
endmodule