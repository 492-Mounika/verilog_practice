// Code your testbench here
// or browse Examples
module tb;
    reg a, b, sel;
    wire z;

    mux_2x1 uut (.a(a), .b(b), .sel(sel), .z(z));

    initial begin
        $monitor("Time=%0t | a=%b b=%b sel=%b => z=%b", $time, a, b, sel, z);

        a = 0; b = 0; sel = 0; #10;
        a = 0; b = 1; sel = 0; #10;
        a = 1; b = 0; sel = 0; #10;
        a = 1; b = 1; sel = 0; #10;

        a = 0; b = 0; sel = 1; #10;
        a = 0; b = 1; sel = 1; #10;
        a = 1; b = 0; sel = 1; #10;
        a = 1; b = 1; sel = 1; #10;

        $finish;
    end
endmodule

  
